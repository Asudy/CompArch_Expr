`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:37:05 08/21/2020 
// Design Name: 
// Module Name:    UnExt 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module UnExt(input [15:0] Imm_16,
				  output[31:0] Imm_32
				 );

	assign Imm_32 = {16'b0, Imm_16};			//��չΪ32λ������
	
endmodule
